//  |---v---|---v---|---v---|---v---|---v---|---v---|---v---|---v---|---v---|---v---|
//-
//-     $_OAI4_ (A, B, C, Y)
//-
//- A 4-input Or-And-Invert gate.
//-
//- Truth table:    A B C D | Y
//-                ---------+---
//-                 0 0 0 0 | 1
//-                 0 0 0 1 | 1
//-                 0 0 1 0 | 1
//-                 0 0 1 1 | 1
//-                 0 1 0 0 | 1
//-                 0 1 0 1 | 0
//-                 0 1 1 0 | 0
//-                 0 1 1 1 | 0
//-                 1 0 0 0 | 1
//-                 1 0 0 1 | 0
//-                 1 0 1 0 | 0
//-                 1 0 1 1 | 0
//-                 1 1 0 0 | 1
//-                 1 1 0 1 | 0
//-                 1 1 1 0 | 0
//-                 1 1 1 1 | 0
//-
module \$_OAI4_ (A, B, C, D, Y);
input A, B, C, D;
output Y;
assign Y = ~((A | B) & (C | D));
endmodule